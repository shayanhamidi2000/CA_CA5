module cacheSim(input[14:0] adr,input clk,rst,output[12:0] HitRate);
    
endmodule
